
module systema (
	button_mode_export,
	clk_clk,
	reset_reset_n,
	btn_op_export);	

	input	[1:0]	button_mode_export;
	input		clk_clk;
	input		reset_reset_n;
	input	[1:0]	btn_op_export;
endmodule
