
module systema (
	button_mode_export,
	clk_clk,
	reset_reset_n);	

	input	[3:0]	button_mode_export;
	input		clk_clk;
	input		reset_reset_n;
endmodule
